module kernel_matrix_trained(conv1_kernel,conv2_kernel,conv3_kernel,connect_matrix);
    parameter bitwidth=32;
    output reg signed [bitwidth-1:0] conv1_kernel [1:0][4:0][4:0];
	output reg signed [bitwidth-1:0] conv2_kernel [1:0][1:0][4:0][4:0];
	output reg signed [bitwidth-1:0] conv3_kernel [9:0][1:0][4:0][4:0];
	output reg signed [bitwidth-1:0] connect_matrix [9:0][9:0];
initial begin
conv1_kernel[0][0][0]=	-73	;
conv1_kernel[0][0][1]=	-51	;
conv1_kernel[0][0][2]=	23	;
conv1_kernel[0][0][3]=	-12	;
conv1_kernel[0][0][4]=	27	;
conv1_kernel[0][1][0]=	-90	;
conv1_kernel[0][1][1]=	24	;
conv1_kernel[0][1][2]=	23	;
conv1_kernel[0][1][3]=	23	;
conv1_kernel[0][1][4]=	13	;
conv1_kernel[0][2][0]=	-71	;
conv1_kernel[0][2][1]=	69	;
conv1_kernel[0][2][2]=	38	;
conv1_kernel[0][2][3]=	37	;
conv1_kernel[0][2][4]=	-5	;
conv1_kernel[0][3][0]=	-27	;
conv1_kernel[0][3][1]=	15	;
conv1_kernel[0][3][2]=	32	;
conv1_kernel[0][3][3]=	17	;
conv1_kernel[0][3][4]=	4	;
conv1_kernel[0][4][0]=	-18	;
conv1_kernel[0][4][1]=	34	;
conv1_kernel[0][4][2]=	-6	;
conv1_kernel[0][4][3]=	-14	;
conv1_kernel[0][4][4]=	-35	;
conv1_kernel[1][0][0]=	14	;
conv1_kernel[1][0][1]=	4	;
conv1_kernel[1][0][2]=	7	;
conv1_kernel[1][0][3]=	-12	;
conv1_kernel[1][0][4]=	-16	;
conv1_kernel[1][1][0]=	26	;
conv1_kernel[1][1][1]=	9	;
conv1_kernel[1][1][2]=	-2	;
conv1_kernel[1][1][3]=	1	;
conv1_kernel[1][1][4]=	-4	;
conv1_kernel[1][2][0]=	23	;
conv1_kernel[1][2][1]=	28	;
conv1_kernel[1][2][2]=	2	;
conv1_kernel[1][2][3]=	0	;
conv1_kernel[1][2][4]=	30	;
conv1_kernel[1][3][0]=	-6	;
conv1_kernel[1][3][1]=	42	;
conv1_kernel[1][3][2]=	67	;
conv1_kernel[1][3][3]=	28	;
conv1_kernel[1][3][4]=	6	;
conv1_kernel[1][4][0]=	0	;
conv1_kernel[1][4][1]=	-6	;
conv1_kernel[1][4][2]=	2	;
conv1_kernel[1][4][3]=	15	;
conv1_kernel[1][4][4]=	15	;
conv2_kernel[0][0][0][0]=	11	;
conv2_kernel[0][0][0][1]=	27	;
conv2_kernel[0][0][0][2]=	34	;
conv2_kernel[0][0][0][3]=	0	;
conv2_kernel[0][0][0][4]=	-3	;
conv2_kernel[0][0][1][0]=	-35	;
conv2_kernel[0][0][1][1]=	25	;
conv2_kernel[0][0][1][2]=	18	;
conv2_kernel[0][0][1][3]=	-11	;
conv2_kernel[0][0][1][4]=	-12	;
conv2_kernel[0][0][2][0]=	8	;
conv2_kernel[0][0][2][1]=	-14	;
conv2_kernel[0][0][2][2]=	-5	;
conv2_kernel[0][0][2][3]=	3	;
conv2_kernel[0][0][2][4]=	22	;
conv2_kernel[0][0][3][0]=	14	;
conv2_kernel[0][0][3][1]=	2	;
conv2_kernel[0][0][3][2]=	-1	;
conv2_kernel[0][0][3][3]=	30	;
conv2_kernel[0][0][3][4]=	11	;
conv2_kernel[0][0][4][0]=	1	;
conv2_kernel[0][0][4][1]=	-30	;
conv2_kernel[0][0][4][2]=	-39	;
conv2_kernel[0][0][4][3]=	-57	;
conv2_kernel[0][0][4][4]=	-8	;
conv2_kernel[0][1][0][0]=	-30	;
conv2_kernel[0][1][0][1]=	-14	;
conv2_kernel[0][1][0][2]=	4	;
conv2_kernel[0][1][0][3]=	16	;
conv2_kernel[0][1][0][4]=	-27	;
conv2_kernel[0][1][1][0]=	-41	;
conv2_kernel[0][1][1][1]=	0	;
conv2_kernel[0][1][1][2]=	3	;
conv2_kernel[0][1][1][3]=	13	;
conv2_kernel[0][1][1][4]=	31	;
conv2_kernel[0][1][2][0]=	32	;
conv2_kernel[0][1][2][1]=	58	;
conv2_kernel[0][1][2][2]=	69	;
conv2_kernel[0][1][2][3]=	79	;
conv2_kernel[0][1][2][4]=	23	;
conv2_kernel[0][1][3][0]=	-18	;
conv2_kernel[0][1][3][1]=	-27	;
conv2_kernel[0][1][3][2]=	-1	;
conv2_kernel[0][1][3][3]=	-30	;
conv2_kernel[0][1][3][4]=	-91	;
conv2_kernel[0][1][4][0]=	-9	;
conv2_kernel[0][1][4][1]=	10	;
conv2_kernel[0][1][4][2]=	-29	;
conv2_kernel[0][1][4][3]=	-45	;
conv2_kernel[0][1][4][4]=	1	;
conv2_kernel[1][0][0][0]=	41	;
conv2_kernel[1][0][0][1]=	28	;
conv2_kernel[1][0][0][2]=	-15	;
conv2_kernel[1][0][0][3]=	-30	;
conv2_kernel[1][0][0][4]=	-12	;
conv2_kernel[1][0][1][0]=	-34	;
conv2_kernel[1][0][1][1]=	-47	;
conv2_kernel[1][0][1][2]=	28	;
conv2_kernel[1][0][1][3]=	-2	;
conv2_kernel[1][0][1][4]=	-29	;
conv2_kernel[1][0][2][0]=	-37	;
conv2_kernel[1][0][2][1]=	-34	;
conv2_kernel[1][0][2][2]=	23	;
conv2_kernel[1][0][2][3]=	24	;
conv2_kernel[1][0][2][4]=	12	;
conv2_kernel[1][0][3][0]=	10	;
conv2_kernel[1][0][3][1]=	-20	;
conv2_kernel[1][0][3][2]=	-62	;
conv2_kernel[1][0][3][3]=	-3	;
conv2_kernel[1][0][3][4]=	4	;
conv2_kernel[1][0][4][0]=	15	;
conv2_kernel[1][0][4][1]=	8	;
conv2_kernel[1][0][4][2]=	6	;
conv2_kernel[1][0][4][3]=	-3	;
conv2_kernel[1][0][4][4]=	4	;
conv2_kernel[1][1][0][0]=	-48	;
conv2_kernel[1][1][0][1]=	-32	;
conv2_kernel[1][1][0][2]=	-41	;
conv2_kernel[1][1][0][3]=	-43	;
conv2_kernel[1][1][0][4]=	-48	;
conv2_kernel[1][1][1][0]=	-12	;
conv2_kernel[1][1][1][1]=	-59	;
conv2_kernel[1][1][1][2]=	10	;
conv2_kernel[1][1][1][3]=	19	;
conv2_kernel[1][1][1][4]=	36	;
conv2_kernel[1][1][2][0]=	124	;
conv2_kernel[1][1][2][1]=	108	;
conv2_kernel[1][1][2][2]=	47	;
conv2_kernel[1][1][2][3]=	5	;
conv2_kernel[1][1][2][4]=	35	;
conv2_kernel[1][1][3][0]=	-50	;
conv2_kernel[1][1][3][1]=	16	;
conv2_kernel[1][1][3][2]=	0	;
conv2_kernel[1][1][3][3]=	15	;
conv2_kernel[1][1][3][4]=	-11	;
conv2_kernel[1][1][4][0]=	-73	;
conv2_kernel[1][1][4][1]=	-13	;
conv2_kernel[1][1][4][2]=	14	;
conv2_kernel[1][1][4][3]=	10	;
conv2_kernel[1][1][4][4]=	-3	;
conv3_kernel[0][0][0][0]=	-65	;
conv3_kernel[0][0][0][1]=	-15	;
conv3_kernel[0][0][0][2]=	19	;
conv3_kernel[0][0][0][3]=	24	;
conv3_kernel[0][0][0][4]=	5	;
conv3_kernel[0][0][1][0]=	-29	;
conv3_kernel[0][0][1][1]=	-3	;
conv3_kernel[0][0][1][2]=	5	;
conv3_kernel[0][0][1][3]=	-7	;
conv3_kernel[0][0][1][4]=	17	;
conv3_kernel[0][0][2][0]=	28	;
conv3_kernel[0][0][2][1]=	17	;
conv3_kernel[0][0][2][2]=	20	;
conv3_kernel[0][0][2][3]=	7	;
conv3_kernel[0][0][2][4]=	1	;
conv3_kernel[0][0][3][0]=	12	;
conv3_kernel[0][0][3][1]=	-5	;
conv3_kernel[0][0][3][2]=	32	;
conv3_kernel[0][0][3][3]=	-23	;
conv3_kernel[0][0][3][4]=	13	;
conv3_kernel[0][0][4][0]=	6	;
conv3_kernel[0][0][4][1]=	-16	;
conv3_kernel[0][0][4][2]=	7	;
conv3_kernel[0][0][4][3]=	2	;
conv3_kernel[0][0][4][4]=	1	;
conv3_kernel[0][1][0][0]=	-19	;
conv3_kernel[0][1][0][1]=	20	;
conv3_kernel[0][1][0][2]=	14	;
conv3_kernel[0][1][0][3]=	-36	;
conv3_kernel[0][1][0][4]=	-17	;
conv3_kernel[0][1][1][0]=	-72	;
conv3_kernel[0][1][1][1]=	6	;
conv3_kernel[0][1][1][2]=	22	;
conv3_kernel[0][1][1][3]=	2	;
conv3_kernel[0][1][1][4]=	-2	;
conv3_kernel[0][1][2][0]=	-48	;
conv3_kernel[0][1][2][1]=	-4	;
conv3_kernel[0][1][2][2]=	27	;
conv3_kernel[0][1][2][3]=	25	;
conv3_kernel[0][1][2][4]=	-47	;
conv3_kernel[0][1][3][0]=	53	;
conv3_kernel[0][1][3][1]=	3	;
conv3_kernel[0][1][3][2]=	-3	;
conv3_kernel[0][1][3][3]=	-17	;
conv3_kernel[0][1][3][4]=	25	;
conv3_kernel[0][1][4][0]=	82	;
conv3_kernel[0][1][4][1]=	-20	;
conv3_kernel[0][1][4][2]=	4	;
conv3_kernel[0][1][4][3]=	13	;
conv3_kernel[0][1][4][4]=	50	;
conv3_kernel[1][0][0][0]=	37	;
conv3_kernel[1][0][0][1]=	19	;
conv3_kernel[1][0][0][2]=	-5	;
conv3_kernel[1][0][0][3]=	-14	;
conv3_kernel[1][0][0][4]=	-83	;
conv3_kernel[1][0][1][0]=	12	;
conv3_kernel[1][0][1][1]=	12	;
conv3_kernel[1][0][1][2]=	-12	;
conv3_kernel[1][0][1][3]=	-4	;
conv3_kernel[1][0][1][4]=	-81	;
conv3_kernel[1][0][2][0]=	-50	;
conv3_kernel[1][0][2][1]=	-11	;
conv3_kernel[1][0][2][2]=	-1	;
conv3_kernel[1][0][2][3]=	2	;
conv3_kernel[1][0][2][4]=	54	;
conv3_kernel[1][0][3][0]=	-25	;
conv3_kernel[1][0][3][1]=	28	;
conv3_kernel[1][0][3][2]=	39	;
conv3_kernel[1][0][3][3]=	-1	;
conv3_kernel[1][0][3][4]=	41	;
conv3_kernel[1][0][4][0]=	39	;
conv3_kernel[1][0][4][1]=	37	;
conv3_kernel[1][0][4][2]=	-8	;
conv3_kernel[1][0][4][3]=	-11	;
conv3_kernel[1][0][4][4]=	-5	;
conv3_kernel[1][1][0][0]=	-26	;
conv3_kernel[1][1][0][1]=	-25	;
conv3_kernel[1][1][0][2]=	-12	;
conv3_kernel[1][1][0][3]=	-7	;
conv3_kernel[1][1][0][4]=	23	;
conv3_kernel[1][1][1][0]=	21	;
conv3_kernel[1][1][1][1]=	-6	;
conv3_kernel[1][1][1][2]=	-20	;
conv3_kernel[1][1][1][3]=	24	;
conv3_kernel[1][1][1][4]=	13	;
conv3_kernel[1][1][2][0]=	25	;
conv3_kernel[1][1][2][1]=	7	;
conv3_kernel[1][1][2][2]=	-14	;
conv3_kernel[1][1][2][3]=	34	;
conv3_kernel[1][1][2][4]=	-16	;
conv3_kernel[1][1][3][0]=	-35	;
conv3_kernel[1][1][3][1]=	26	;
conv3_kernel[1][1][3][2]=	-12	;
conv3_kernel[1][1][3][3]=	-6	;
conv3_kernel[1][1][3][4]=	16	;
conv3_kernel[1][1][4][0]=	-90	;
conv3_kernel[1][1][4][1]=	21	;
conv3_kernel[1][1][4][2]=	14	;
conv3_kernel[1][1][4][3]=	43	;
conv3_kernel[1][1][4][4]=	39	;
conv3_kernel[2][0][0][0]=	30	;
conv3_kernel[2][0][0][1]=	42	;
conv3_kernel[2][0][0][2]=	-16	;
conv3_kernel[2][0][0][3]=	18	;
conv3_kernel[2][0][0][4]=	-37	;
conv3_kernel[2][0][1][0]=	-16	;
conv3_kernel[2][0][1][1]=	14	;
conv3_kernel[2][0][1][2]=	10	;
conv3_kernel[2][0][1][3]=	-3	;
conv3_kernel[2][0][1][4]=	-43	;
conv3_kernel[2][0][2][0]=	7	;
conv3_kernel[2][0][2][1]=	7	;
conv3_kernel[2][0][2][2]=	-11	;
conv3_kernel[2][0][2][3]=	59	;
conv3_kernel[2][0][2][4]=	35	;
conv3_kernel[2][0][3][0]=	9	;
conv3_kernel[2][0][3][1]=	-2	;
conv3_kernel[2][0][3][2]=	2	;
conv3_kernel[2][0][3][3]=	59	;
conv3_kernel[2][0][3][4]=	17	;
conv3_kernel[2][0][4][0]=	-6	;
conv3_kernel[2][0][4][1]=	-22	;
conv3_kernel[2][0][4][2]=	-30	;
conv3_kernel[2][0][4][3]=	-4	;
conv3_kernel[2][0][4][4]=	15	;
conv3_kernel[2][1][0][0]=	-2	;
conv3_kernel[2][1][0][1]=	0	;
conv3_kernel[2][1][0][2]=	8	;
conv3_kernel[2][1][0][3]=	0	;
conv3_kernel[2][1][0][4]=	15	;
conv3_kernel[2][1][1][0]=	29	;
conv3_kernel[2][1][1][1]=	10	;
conv3_kernel[2][1][1][2]=	11	;
conv3_kernel[2][1][1][3]=	29	;
conv3_kernel[2][1][1][4]=	10	;
conv3_kernel[2][1][2][0]=	-24	;
conv3_kernel[2][1][2][1]=	-6	;
conv3_kernel[2][1][2][2]=	9	;
conv3_kernel[2][1][2][3]=	47	;
conv3_kernel[2][1][2][4]=	-45	;
conv3_kernel[2][1][3][0]=	-7	;
conv3_kernel[2][1][3][1]=	7	;
conv3_kernel[2][1][3][2]=	15	;
conv3_kernel[2][1][3][3]=	-30	;
conv3_kernel[2][1][3][4]=	-35	;
conv3_kernel[2][1][4][0]=	25	;
conv3_kernel[2][1][4][1]=	-16	;
conv3_kernel[2][1][4][2]=	-34	;
conv3_kernel[2][1][4][3]=	-7	;
conv3_kernel[2][1][4][4]=	-1	;
conv3_kernel[3][0][0][0]=	10	;
conv3_kernel[3][0][0][1]=	-16	;
conv3_kernel[3][0][0][2]=	13	;
conv3_kernel[3][0][0][3]=	-13	;
conv3_kernel[3][0][0][4]=	-20	;
conv3_kernel[3][0][1][0]=	22	;
conv3_kernel[3][0][1][1]=	-11	;
conv3_kernel[3][0][1][2]=	0	;
conv3_kernel[3][0][1][3]=	1	;
conv3_kernel[3][0][1][4]=	34	;
conv3_kernel[3][0][2][0]=	-1	;
conv3_kernel[3][0][2][1]=	-32	;
conv3_kernel[3][0][2][2]=	1	;
conv3_kernel[3][0][2][3]=	26	;
conv3_kernel[3][0][2][4]=	17	;
conv3_kernel[3][0][3][0]=	-20	;
conv3_kernel[3][0][3][1]=	-9	;
conv3_kernel[3][0][3][2]=	16	;
conv3_kernel[3][0][3][3]=	-58	;
conv3_kernel[3][0][3][4]=	-9	;
conv3_kernel[3][0][4][0]=	33	;
conv3_kernel[3][0][4][1]=	19	;
conv3_kernel[3][0][4][2]=	29	;
conv3_kernel[3][0][4][3]=	-7	;
conv3_kernel[3][0][4][4]=	-32	;
conv3_kernel[3][1][0][0]=	17	;
conv3_kernel[3][1][0][1]=	8	;
conv3_kernel[3][1][0][2]=	8	;
conv3_kernel[3][1][0][3]=	-40	;
conv3_kernel[3][1][0][4]=	17	;
conv3_kernel[3][1][1][0]=	-13	;
conv3_kernel[3][1][1][1]=	2	;
conv3_kernel[3][1][1][2]=	16	;
conv3_kernel[3][1][1][3]=	12	;
conv3_kernel[3][1][1][4]=	-6	;
conv3_kernel[3][1][2][0]=	-16	;
conv3_kernel[3][1][2][1]=	0	;
conv3_kernel[3][1][2][2]=	59	;
conv3_kernel[3][1][2][3]=	42	;
conv3_kernel[3][1][2][4]=	29	;
conv3_kernel[3][1][3][0]=	66	;
conv3_kernel[3][1][3][1]=	-8	;
conv3_kernel[3][1][3][2]=	-9	;
conv3_kernel[3][1][3][3]=	19	;
conv3_kernel[3][1][3][4]=	55	;
conv3_kernel[3][1][4][0]=	-121	;
conv3_kernel[3][1][4][1]=	-13	;
conv3_kernel[3][1][4][2]=	11	;
conv3_kernel[3][1][4][3]=	12	;
conv3_kernel[3][1][4][4]=	-12	;
conv3_kernel[4][0][0][0]=	-8	;
conv3_kernel[4][0][0][1]=	32	;
conv3_kernel[4][0][0][2]=	50	;
conv3_kernel[4][0][0][3]=	78	;
conv3_kernel[4][0][0][4]=	50	;
conv3_kernel[4][0][1][0]=	10	;
conv3_kernel[4][0][1][1]=	4	;
conv3_kernel[4][0][1][2]=	5	;
conv3_kernel[4][0][1][3]=	11	;
conv3_kernel[4][0][1][4]=	24	;
conv3_kernel[4][0][2][0]=	-25	;
conv3_kernel[4][0][2][1]=	-8	;
conv3_kernel[4][0][2][2]=	22	;
conv3_kernel[4][0][2][3]=	-36	;
conv3_kernel[4][0][2][4]=	-45	;
conv3_kernel[4][0][3][0]=	-10	;
conv3_kernel[4][0][3][1]=	1	;
conv3_kernel[4][0][3][2]=	37	;
conv3_kernel[4][0][3][3]=	-24	;
conv3_kernel[4][0][3][4]=	-1	;
conv3_kernel[4][0][4][0]=	9	;
conv3_kernel[4][0][4][1]=	-11	;
conv3_kernel[4][0][4][2]=	20	;
conv3_kernel[4][0][4][3]=	5	;
conv3_kernel[4][0][4][4]=	-29	;
conv3_kernel[4][1][0][0]=	22	;
conv3_kernel[4][1][0][1]=	-15	;
conv3_kernel[4][1][0][2]=	-34	;
conv3_kernel[4][1][0][3]=	-75	;
conv3_kernel[4][1][0][4]=	-18	;
conv3_kernel[4][1][1][0]=	-21	;
conv3_kernel[4][1][1][1]=	-13	;
conv3_kernel[4][1][1][2]=	-7	;
conv3_kernel[4][1][1][3]=	14	;
conv3_kernel[4][1][1][4]=	73	;
conv3_kernel[4][1][2][0]=	-37	;
conv3_kernel[4][1][2][1]=	6	;
conv3_kernel[4][1][2][2]=	31	;
conv3_kernel[4][1][2][3]=	50	;
conv3_kernel[4][1][2][4]=	48	;
conv3_kernel[4][1][3][0]=	-3	;
conv3_kernel[4][1][3][1]=	33	;
conv3_kernel[4][1][3][2]=	5	;
conv3_kernel[4][1][3][3]=	18	;
conv3_kernel[4][1][3][4]=	-10	;
conv3_kernel[4][1][4][0]=	-35	;
conv3_kernel[4][1][4][1]=	23	;
conv3_kernel[4][1][4][2]=	12	;
conv3_kernel[4][1][4][3]=	26	;
conv3_kernel[4][1][4][4]=	-3	;
conv3_kernel[5][0][0][0]=	77	;
conv3_kernel[5][0][0][1]=	33	;
conv3_kernel[5][0][0][2]=	23	;
conv3_kernel[5][0][0][3]=	-17	;
conv3_kernel[5][0][0][4]=	-34	;
conv3_kernel[5][0][1][0]=	45	;
conv3_kernel[5][0][1][1]=	12	;
conv3_kernel[5][0][1][2]=	4	;
conv3_kernel[5][0][1][3]=	-3	;
conv3_kernel[5][0][1][4]=	8	;
conv3_kernel[5][0][2][0]=	15	;
conv3_kernel[5][0][2][1]=	-6	;
conv3_kernel[5][0][2][2]=	-9	;
conv3_kernel[5][0][2][3]=	3	;
conv3_kernel[5][0][2][4]=	-22	;
conv3_kernel[5][0][3][0]=	0	;
conv3_kernel[5][0][3][1]=	13	;
conv3_kernel[5][0][3][2]=	-9	;
conv3_kernel[5][0][3][3]=	-3	;
conv3_kernel[5][0][3][4]=	-2	;
conv3_kernel[5][0][4][0]=	3	;
conv3_kernel[5][0][4][1]=	-23	;
conv3_kernel[5][0][4][2]=	-23	;
conv3_kernel[5][0][4][3]=	8	;
conv3_kernel[5][0][4][4]=	-34	;
conv3_kernel[5][1][0][0]=	-44	;
conv3_kernel[5][1][0][1]=	5	;
conv3_kernel[5][1][0][2]=	16	;
conv3_kernel[5][1][0][3]=	-3	;
conv3_kernel[5][1][0][4]=	6	;
conv3_kernel[5][1][1][0]=	-18	;
conv3_kernel[5][1][1][1]=	31	;
conv3_kernel[5][1][1][2]=	12	;
conv3_kernel[5][1][1][3]=	21	;
conv3_kernel[5][1][1][4]=	9	;
conv3_kernel[5][1][2][0]=	61	;
conv3_kernel[5][1][2][1]=	-7	;
conv3_kernel[5][1][2][2]=	2	;
conv3_kernel[5][1][2][3]=	18	;
conv3_kernel[5][1][2][4]=	37	;
conv3_kernel[5][1][3][0]=	96	;
conv3_kernel[5][1][3][1]=	12	;
conv3_kernel[5][1][3][2]=	-13	;
conv3_kernel[5][1][3][3]=	24	;
conv3_kernel[5][1][3][4]=	10	;
conv3_kernel[5][1][4][0]=	84	;
conv3_kernel[5][1][4][1]=	25	;
conv3_kernel[5][1][4][2]=	19	;
conv3_kernel[5][1][4][3]=	2	;
conv3_kernel[5][1][4][4]=	-21	;
conv3_kernel[6][0][0][0]=	-11	;
conv3_kernel[6][0][0][1]=	-47	;
conv3_kernel[6][0][0][2]=	-24	;
conv3_kernel[6][0][0][3]=	6	;
conv3_kernel[6][0][0][4]=	35	;
conv3_kernel[6][0][1][0]=	-15	;
conv3_kernel[6][0][1][1]=	17	;
conv3_kernel[6][0][1][2]=	9	;
conv3_kernel[6][0][1][3]=	9	;
conv3_kernel[6][0][1][4]=	23	;
conv3_kernel[6][0][2][0]=	17	;
conv3_kernel[6][0][2][1]=	-2	;
conv3_kernel[6][0][2][2]=	-14	;
conv3_kernel[6][0][2][3]=	58	;
conv3_kernel[6][0][2][4]=	18	;
conv3_kernel[6][0][3][0]=	-8	;
conv3_kernel[6][0][3][1]=	18	;
conv3_kernel[6][0][3][2]=	-6	;
conv3_kernel[6][0][3][3]=	24	;
conv3_kernel[6][0][3][4]=	38	;
conv3_kernel[6][0][4][0]=	30	;
conv3_kernel[6][0][4][1]=	-11	;
conv3_kernel[6][0][4][2]=	0	;
conv3_kernel[6][0][4][3]=	9	;
conv3_kernel[6][0][4][4]=	-9	;
conv3_kernel[6][1][0][0]=	44	;
conv3_kernel[6][1][0][1]=	8	;
conv3_kernel[6][1][0][2]=	-31	;
conv3_kernel[6][1][0][3]=	-72	;
conv3_kernel[6][1][0][4]=	-37	;
conv3_kernel[6][1][1][0]=	-20	;
conv3_kernel[6][1][1][1]=	2	;
conv3_kernel[6][1][1][2]=	-6	;
conv3_kernel[6][1][1][3]=	-11	;
conv3_kernel[6][1][1][4]=	-9	;
conv3_kernel[6][1][2][0]=	39	;
conv3_kernel[6][1][2][1]=	13	;
conv3_kernel[6][1][2][2]=	18	;
conv3_kernel[6][1][2][3]=	68	;
conv3_kernel[6][1][2][4]=	10	;
conv3_kernel[6][1][3][0]=	45	;
conv3_kernel[6][1][3][1]=	15	;
conv3_kernel[6][1][3][2]=	9	;
conv3_kernel[6][1][3][3]=	22	;
conv3_kernel[6][1][3][4]=	49	;
conv3_kernel[6][1][4][0]=	-31	;
conv3_kernel[6][1][4][1]=	-15	;
conv3_kernel[6][1][4][2]=	-11	;
conv3_kernel[6][1][4][3]=	-39	;
conv3_kernel[6][1][4][4]=	22	;
conv3_kernel[7][0][0][0]=	-15	;
conv3_kernel[7][0][0][1]=	-1	;
conv3_kernel[7][0][0][2]=	-41	;
conv3_kernel[7][0][0][3]=	-22	;
conv3_kernel[7][0][0][4]=	-4	;
conv3_kernel[7][0][1][0]=	-71	;
conv3_kernel[7][0][1][1]=	4	;
conv3_kernel[7][0][1][2]=	18	;
conv3_kernel[7][0][1][3]=	9	;
conv3_kernel[7][0][1][4]=	4	;
conv3_kernel[7][0][2][0]=	13	;
conv3_kernel[7][0][2][1]=	12	;
conv3_kernel[7][0][2][2]=	9	;
conv3_kernel[7][0][2][3]=	7	;
conv3_kernel[7][0][2][4]=	16	;
conv3_kernel[7][0][3][0]=	25	;
conv3_kernel[7][0][3][1]=	3	;
conv3_kernel[7][0][3][2]=	-2	;
conv3_kernel[7][0][3][3]=	-23	;
conv3_kernel[7][0][3][4]=	-62	;
conv3_kernel[7][0][4][0]=	-2	;
conv3_kernel[7][0][4][1]=	2	;
conv3_kernel[7][0][4][2]=	-14	;
conv3_kernel[7][0][4][3]=	6	;
conv3_kernel[7][0][4][4]=	33	;
conv3_kernel[7][1][0][0]=	10	;
conv3_kernel[7][1][0][1]=	40	;
conv3_kernel[7][1][0][2]=	5	;
conv3_kernel[7][1][0][3]=	2	;
conv3_kernel[7][1][0][4]=	35	;
conv3_kernel[7][1][1][0]=	39	;
conv3_kernel[7][1][1][1]=	5	;
conv3_kernel[7][1][1][2]=	8	;
conv3_kernel[7][1][1][3]=	9	;
conv3_kernel[7][1][1][4]=	15	;
conv3_kernel[7][1][2][0]=	-37	;
conv3_kernel[7][1][2][1]=	-27	;
conv3_kernel[7][1][2][2]=	34	;
conv3_kernel[7][1][2][3]=	56	;
conv3_kernel[7][1][2][4]=	-6	;
conv3_kernel[7][1][3][0]=	-23	;
conv3_kernel[7][1][3][1]=	24	;
conv3_kernel[7][1][3][2]=	35	;
conv3_kernel[7][1][3][3]=	21	;
conv3_kernel[7][1][3][4]=	-42	;
conv3_kernel[7][1][4][0]=	37	;
conv3_kernel[7][1][4][1]=	20	;
conv3_kernel[7][1][4][2]=	27	;
conv3_kernel[7][1][4][3]=	-10	;
conv3_kernel[7][1][4][4]=	-70	;
conv3_kernel[8][0][0][0]=	-76	;
conv3_kernel[8][0][0][1]=	-29	;
conv3_kernel[8][0][0][2]=	15	;
conv3_kernel[8][0][0][3]=	-3	;
conv3_kernel[8][0][0][4]=	22	;
conv3_kernel[8][0][1][0]=	-116	;
conv3_kernel[8][0][1][1]=	2	;
conv3_kernel[8][0][1][2]=	2	;
conv3_kernel[8][0][1][3]=	5	;
conv3_kernel[8][0][1][4]=	-8	;
conv3_kernel[8][0][2][0]=	22	;
conv3_kernel[8][0][2][1]=	-18	;
conv3_kernel[8][0][2][2]=	16	;
conv3_kernel[8][0][2][3]=	13	;
conv3_kernel[8][0][2][4]=	40	;
conv3_kernel[8][0][3][0]=	-2	;
conv3_kernel[8][0][3][1]=	-3	;
conv3_kernel[8][0][3][2]=	10	;
conv3_kernel[8][0][3][3]=	-15	;
conv3_kernel[8][0][3][4]=	-3	;
conv3_kernel[8][0][4][0]=	18	;
conv3_kernel[8][0][4][1]=	7	;
conv3_kernel[8][0][4][2]=	-2	;
conv3_kernel[8][0][4][3]=	8	;
conv3_kernel[8][0][4][4]=	-5	;
conv3_kernel[8][1][0][0]=	57	;
conv3_kernel[8][1][0][1]=	40	;
conv3_kernel[8][1][0][2]=	3	;
conv3_kernel[8][1][0][3]=	-6	;
conv3_kernel[8][1][0][4]=	30	;
conv3_kernel[8][1][1][0]=	25	;
conv3_kernel[8][1][1][1]=	7	;
conv3_kernel[8][1][1][2]=	10	;
conv3_kernel[8][1][1][3]=	27	;
conv3_kernel[8][1][1][4]=	31	;
conv3_kernel[8][1][2][0]=	6	;
conv3_kernel[8][1][2][1]=	-33	;
conv3_kernel[8][1][2][2]=	-40	;
conv3_kernel[8][1][2][3]=	-16	;
conv3_kernel[8][1][2][4]=	-32	;
conv3_kernel[8][1][3][0]=	-17	;
conv3_kernel[8][1][3][1]=	-14	;
conv3_kernel[8][1][3][2]=	-16	;
conv3_kernel[8][1][3][3]=	0	;
conv3_kernel[8][1][3][4]=	-27	;
conv3_kernel[8][1][4][0]=	-76	;
conv3_kernel[8][1][4][1]=	9	;
conv3_kernel[8][1][4][2]=	9	;
conv3_kernel[8][1][4][3]=	11	;
conv3_kernel[8][1][4][4]=	-60	;
conv3_kernel[9][0][0][0]=	43	;
conv3_kernel[9][0][0][1]=	-28	;
conv3_kernel[9][0][0][2]=	-28	;
conv3_kernel[9][0][0][3]=	-49	;
conv3_kernel[9][0][0][4]=	-24	;
conv3_kernel[9][0][1][0]=	41	;
conv3_kernel[9][0][1][1]=	-18	;
conv3_kernel[9][0][1][2]=	17	;
conv3_kernel[9][0][1][3]=	18	;
conv3_kernel[9][0][1][4]=	9	;
conv3_kernel[9][0][2][0]=	-3	;
conv3_kernel[9][0][2][1]=	-14	;
conv3_kernel[9][0][2][2]=	70	;
conv3_kernel[9][0][2][3]=	41	;
conv3_kernel[9][0][2][4]=	0	;
conv3_kernel[9][0][3][0]=	-19	;
conv3_kernel[9][0][3][1]=	-16	;
conv3_kernel[9][0][3][2]=	42	;
conv3_kernel[9][0][3][3]=	-30	;
conv3_kernel[9][0][3][4]=	1	;
conv3_kernel[9][0][4][0]=	4	;
conv3_kernel[9][0][4][1]=	-38	;
conv3_kernel[9][0][4][2]=	44	;
conv3_kernel[9][0][4][3]=	24	;
conv3_kernel[9][0][4][4]=	-22	;
conv3_kernel[9][1][0][0]=	-7	;
conv3_kernel[9][1][0][1]=	13	;
conv3_kernel[9][1][0][2]=	44	;
conv3_kernel[9][1][0][3]=	-36	;
conv3_kernel[9][1][0][4]=	-8	;
conv3_kernel[9][1][1][0]=	-5	;
conv3_kernel[9][1][1][1]=	-12	;
conv3_kernel[9][1][1][2]=	11	;
conv3_kernel[9][1][1][3]=	-25	;
conv3_kernel[9][1][1][4]=	-35	;
conv3_kernel[9][1][2][0]=	-2	;
conv3_kernel[9][1][2][1]=	-12	;
conv3_kernel[9][1][2][2]=	29	;
conv3_kernel[9][1][2][3]=	-3	;
conv3_kernel[9][1][2][4]=	-1	;
conv3_kernel[9][1][3][0]=	17	;
conv3_kernel[9][1][3][1]=	7	;
conv3_kernel[9][1][3][2]=	4	;
conv3_kernel[9][1][3][3]=	4	;
conv3_kernel[9][1][3][4]=	3	;
conv3_kernel[9][1][4][0]=	14	;
conv3_kernel[9][1][4][1]=	27	;
conv3_kernel[9][1][4][2]=	1	;
conv3_kernel[9][1][4][3]=	-4	;
conv3_kernel[9][1][4][4]=	-13	;
connect_matrix [0][0]=	-43	;
connect_matrix [0][1]=	49	;
connect_matrix [0][2]=	-7	;
connect_matrix [0][3]=	-39	;
connect_matrix [0][4]=	7	;
connect_matrix [0][5]=	-8	;
connect_matrix [0][6]=	-3	;
connect_matrix [0][7]=	-2	;
connect_matrix [0][8]=	25	;
connect_matrix [0][9]=	-24	;
connect_matrix [1][0]=	54	;
connect_matrix [1][1]=	-18	;
connect_matrix [1][2]=	-51	;
connect_matrix [1][3]=	-39	;
connect_matrix [1][4]=	0	;
connect_matrix [1][5]=	19	;
connect_matrix [1][6]=	20	;
connect_matrix [1][7]=	-94	;
connect_matrix [1][8]=	50	;
connect_matrix [1][9]=	74	;
connect_matrix [2][0]=	20	;
connect_matrix [2][1]=	42	;
connect_matrix [2][2]=	-2	;
connect_matrix [2][3]=	19	;
connect_matrix [2][4]=	-45	;
connect_matrix [2][5]=	24	;
connect_matrix [2][6]=	6	;
connect_matrix [2][7]=	-22	;
connect_matrix [2][8]=	-57	;
connect_matrix [2][9]=	-3	;
connect_matrix [3][0]=	-14	;
connect_matrix [3][1]=	-2	;
connect_matrix [3][2]=	-32	;
connect_matrix [3][3]=	-1	;
connect_matrix [3][4]=	-9	;
connect_matrix [3][5]=	47	;
connect_matrix [3][6]=	-13	;
connect_matrix [3][7]=	22	;
connect_matrix [3][8]=	-45	;
connect_matrix [3][9]=	22	;
connect_matrix [4][0]=	0	;
connect_matrix [4][1]=	-18	;
connect_matrix [4][2]=	-5	;
connect_matrix [4][3]=	-17	;
connect_matrix [4][4]=	-34	;
connect_matrix [4][5]=	-46	;
connect_matrix [4][6]=	64	;
connect_matrix [4][7]=	28	;
connect_matrix [4][8]=	-20	;
connect_matrix [4][9]=	23	;
connect_matrix [5][0]=	18	;
connect_matrix [5][1]=	-32	;
connect_matrix [5][2]=	-34	;
connect_matrix [5][3]=	-13	;
connect_matrix [5][4]=	42	;
connect_matrix [5][5]=	25	;
connect_matrix [5][6]=	-7	;
connect_matrix [5][7]=	20	;
connect_matrix [5][8]=	-6	;
connect_matrix [5][9]=	-38	;
connect_matrix [6][0]=	-52	;
connect_matrix [6][1]=	26	;
connect_matrix [6][2]=	21	;
connect_matrix [6][3]=	9	;
connect_matrix [6][4]=	62	;
connect_matrix [6][5]=	-91	;
connect_matrix [6][6]=	13	;
connect_matrix [6][7]=	-14	;
connect_matrix [6][8]=	-14	;
connect_matrix [6][9]=	-16	;
connect_matrix [7][0]=	-32	;
connect_matrix [7][1]=	-43	;
connect_matrix [7][2]=	54	;
connect_matrix [7][3]=	20	;
connect_matrix [7][4]=	-5	;
connect_matrix [7][5]=	28	;
connect_matrix [7][6]=	0	;
connect_matrix [7][7]=	-39	;
connect_matrix [7][8]=	27	;
connect_matrix [7][9]=	17	;
connect_matrix [8][0]=	7	;
connect_matrix [8][1]=	-2	;
connect_matrix [8][2]=	2	;
connect_matrix [8][3]=	58	;
connect_matrix [8][4]=	-14	;
connect_matrix [8][5]=	-9	;
connect_matrix [8][6]=	-29	;
connect_matrix [8][7]=	12	;
connect_matrix [8][8]=	11	;
connect_matrix [8][9]=	-9	;
connect_matrix [9][0]=	27	;
connect_matrix [9][1]=	-7	;
connect_matrix [9][2]=	38	;
connect_matrix [9][3]=	-20	;
connect_matrix [9][4]=	-11	;
connect_matrix [9][5]=	-23	;
connect_matrix [9][6]=	-35	;
connect_matrix [9][7]=	42	;
connect_matrix [9][8]=	-31	;
connect_matrix [9][9]=	17	;

end
endmodule