module kernel_matrix_trained(conv1_kernel,conv2_kernel,conv3_kernel,connect_matrix);
parameter bitwidth=32;
output reg signed [bitwidth-1:0] conv1_kernel [1:0][4:0][4:0];
output reg signed [bitwidth-1:0] conv2_kernel [1:0][1:0][4:0][4:0];
output reg signed [bitwidth-1:0] conv3_kernel [9:0][1:0][4:0][4:0];
output reg signed [bitwidth-1:0] connect_matrix [9:0][9:0];
//always@(*) begin
initial begin
conv1_kernel[0][0][0]=	-9357	;
conv1_kernel[0][0][1]=	-6475	;
conv1_kernel[0][0][2]=	2935	;
conv1_kernel[0][0][3]=	-1600	;
conv1_kernel[0][0][4]=	3413	;
conv1_kernel[0][1][0]=	-11490	;
conv1_kernel[0][1][1]=	3066	;
conv1_kernel[0][1][2]=	2881	;
conv1_kernel[0][1][3]=	2993	;
conv1_kernel[0][1][4]=	1627	;
conv1_kernel[0][2][0]=	-9081	;
conv1_kernel[0][2][1]=	8797	;
conv1_kernel[0][2][2]=	4886	;
conv1_kernel[0][2][3]=	4693	;
conv1_kernel[0][2][4]=	-625	;
conv1_kernel[0][3][0]=	-3471	;
conv1_kernel[0][3][1]=	1973	;
conv1_kernel[0][3][2]=	4050	;
conv1_kernel[0][3][3]=	2125	;
conv1_kernel[0][3][4]=	567	;
conv1_kernel[0][4][0]=	-2259	;
conv1_kernel[0][4][1]=	4348	;
conv1_kernel[0][4][2]=	-826	;
conv1_kernel[0][4][3]=	-1821	;
conv1_kernel[0][4][4]=	-4515	;
conv1_kernel[1][0][0]=	1789	;
conv1_kernel[1][0][1]=	570	;
conv1_kernel[1][0][2]=	869	;
conv1_kernel[1][0][3]=	-1511	;
conv1_kernel[1][0][4]=	-2055	;
conv1_kernel[1][1][0]=	3382	;
conv1_kernel[1][1][1]=	1134	;
conv1_kernel[1][1][2]=	-244	;
conv1_kernel[1][1][3]=	69	;
conv1_kernel[1][1][4]=	-482	;
conv1_kernel[1][2][0]=	2973	;
conv1_kernel[1][2][1]=	3625	;
conv1_kernel[1][2][2]=	275	;
conv1_kernel[1][2][3]=	60	;
conv1_kernel[1][2][4]=	3885	;
conv1_kernel[1][3][0]=	-798	;
conv1_kernel[1][3][1]=	5364	;
conv1_kernel[1][3][2]=	8564	;
conv1_kernel[1][3][3]=	3612	;
conv1_kernel[1][3][4]=	808	;
conv1_kernel[1][4][0]=	-32	;
conv1_kernel[1][4][1]=	-735	;
conv1_kernel[1][4][2]=	256	;
conv1_kernel[1][4][3]=	1911	;
conv1_kernel[1][4][4]=	1983	;
conv2_kernel[0][0][0][0]=	1420	;
conv2_kernel[0][0][0][1]=	3444	;
conv2_kernel[0][0][0][2]=	4399	;
conv2_kernel[0][0][0][3]=	-14	;
conv2_kernel[0][0][0][4]=	-383	;
conv2_kernel[0][0][1][0]=	-4492	;
conv2_kernel[0][0][1][1]=	3191	;
conv2_kernel[0][0][1][2]=	2244	;
conv2_kernel[0][0][1][3]=	-1452	;
conv2_kernel[0][0][1][4]=	-1506	;
conv2_kernel[0][0][2][0]=	1025	;
conv2_kernel[0][0][2][1]=	-1853	;
conv2_kernel[0][0][2][2]=	-631	;
conv2_kernel[0][0][2][3]=	408	;
conv2_kernel[0][0][2][4]=	2873	;
conv2_kernel[0][0][3][0]=	1776	;
conv2_kernel[0][0][3][1]=	310	;
conv2_kernel[0][0][3][2]=	-71	;
conv2_kernel[0][0][3][3]=	3814	;
conv2_kernel[0][0][3][4]=	1400	;
conv2_kernel[0][0][4][0]=	159	;
conv2_kernel[0][0][4][1]=	-3865	;
conv2_kernel[0][0][4][2]=	-5031	;
conv2_kernel[0][0][4][3]=	-7287	;
conv2_kernel[0][0][4][4]=	-1074	;
conv2_kernel[0][1][0][0]=	-3879	;
conv2_kernel[0][1][0][1]=	-1853	;
conv2_kernel[0][1][0][2]=	508	;
conv2_kernel[0][1][0][3]=	2066	;
conv2_kernel[0][1][0][4]=	-3506	;
conv2_kernel[0][1][1][0]=	-5217	;
conv2_kernel[0][1][1][1]=	3	;
conv2_kernel[0][1][1][2]=	398	;
conv2_kernel[0][1][1][3]=	1692	;
conv2_kernel[0][1][1][4]=	3957	;
conv2_kernel[0][1][2][0]=	4042	;
conv2_kernel[0][1][2][1]=	7483	;
conv2_kernel[0][1][2][2]=	8781	;
conv2_kernel[0][1][2][3]=	10138	;
conv2_kernel[0][1][2][4]=	2943	;
conv2_kernel[0][1][3][0]=	-2276	;
conv2_kernel[0][1][3][1]=	-3427	;
conv2_kernel[0][1][3][2]=	-93	;
conv2_kernel[0][1][3][3]=	-3834	;
conv2_kernel[0][1][3][4]=	-11595	;
conv2_kernel[0][1][4][0]=	-1106	;
conv2_kernel[0][1][4][1]=	1218	;
conv2_kernel[0][1][4][2]=	-3736	;
conv2_kernel[0][1][4][3]=	-5789	;
conv2_kernel[0][1][4][4]=	181	;
conv2_kernel[1][0][0][0]=	5184	;
conv2_kernel[1][0][0][1]=	3569	;
conv2_kernel[1][0][0][2]=	-1898	;
conv2_kernel[1][0][0][3]=	-3864	;
conv2_kernel[1][0][0][4]=	-1522	;
conv2_kernel[1][0][1][0]=	-4330	;
conv2_kernel[1][0][1][1]=	-5999	;
conv2_kernel[1][0][1][2]=	3530	;
conv2_kernel[1][0][1][3]=	-281	;
conv2_kernel[1][0][1][4]=	-3691	;
conv2_kernel[1][0][2][0]=	-4780	;
conv2_kernel[1][0][2][1]=	-4325	;
conv2_kernel[1][0][2][2]=	2948	;
conv2_kernel[1][0][2][3]=	3135	;
conv2_kernel[1][0][2][4]=	1481	;
conv2_kernel[1][0][3][0]=	1223	;
conv2_kernel[1][0][3][1]=	-2568	;
conv2_kernel[1][0][3][2]=	-7893	;
conv2_kernel[1][0][3][3]=	-442	;
conv2_kernel[1][0][3][4]=	519	;
conv2_kernel[1][0][4][0]=	1944	;
conv2_kernel[1][0][4][1]=	1057	;
conv2_kernel[1][0][4][2]=	781	;
conv2_kernel[1][0][4][3]=	-335	;
conv2_kernel[1][0][4][4]=	472	;
conv2_kernel[1][1][0][0]=	-6090	;
conv2_kernel[1][1][0][1]=	-4126	;
conv2_kernel[1][1][0][2]=	-5310	;
conv2_kernel[1][1][0][3]=	-5478	;
conv2_kernel[1][1][0][4]=	-6192	;
conv2_kernel[1][1][1][0]=	-1492	;
conv2_kernel[1][1][1][1]=	-7515	;
conv2_kernel[1][1][1][2]=	1326	;
conv2_kernel[1][1][1][3]=	2419	;
conv2_kernel[1][1][1][4]=	4545	;
conv2_kernel[1][1][2][0]=	15903	;
conv2_kernel[1][1][2][1]=	13792	;
conv2_kernel[1][1][2][2]=	6033	;
conv2_kernel[1][1][2][3]=	613	;
conv2_kernel[1][1][2][4]=	4478	;
conv2_kernel[1][1][3][0]=	-6364	;
conv2_kernel[1][1][3][1]=	2088	;
conv2_kernel[1][1][3][2]=	16	;
conv2_kernel[1][1][3][3]=	1878	;
conv2_kernel[1][1][3][4]=	-1416	;
conv2_kernel[1][1][4][0]=	-9317	;
conv2_kernel[1][1][4][1]=	-1645	;
conv2_kernel[1][1][4][2]=	1790	;
conv2_kernel[1][1][4][3]=	1292	;
conv2_kernel[1][1][4][4]=	-431	;
conv3_kernel[0][0][0][0]=	-8372	;
conv3_kernel[0][0][0][1]=	-1915	;
conv3_kernel[0][0][0][2]=	2435	;
conv3_kernel[0][0][0][3]=	3130	;
conv3_kernel[0][0][0][4]=	703	;
conv3_kernel[0][0][1][0]=	-3714	;
conv3_kernel[0][0][1][1]=	-399	;
conv3_kernel[0][0][1][2]=	633	;
conv3_kernel[0][0][1][3]=	-841	;
conv3_kernel[0][0][1][4]=	2236	;
conv3_kernel[0][0][2][0]=	3556	;
conv3_kernel[0][0][2][1]=	2216	;
conv3_kernel[0][0][2][2]=	2538	;
conv3_kernel[0][0][2][3]=	927	;
conv3_kernel[0][0][2][4]=	145	;
conv3_kernel[0][0][3][0]=	1575	;
conv3_kernel[0][0][3][1]=	-585	;
conv3_kernel[0][0][3][2]=	4042	;
conv3_kernel[0][0][3][3]=	-2882	;
conv3_kernel[0][0][3][4]=	1717	;
conv3_kernel[0][0][4][0]=	830	;
conv3_kernel[0][0][4][1]=	-2065	;
conv3_kernel[0][0][4][2]=	919	;
conv3_kernel[0][0][4][3]=	231	;
conv3_kernel[0][0][4][4]=	165	;
conv3_kernel[0][1][0][0]=	-2462	;
conv3_kernel[0][1][0][1]=	2550	;
conv3_kernel[0][1][0][2]=	1767	;
conv3_kernel[0][1][0][3]=	-4544	;
conv3_kernel[0][1][0][4]=	-2225	;
conv3_kernel[0][1][1][0]=	-9195	;
conv3_kernel[0][1][1][1]=	746	;
conv3_kernel[0][1][1][2]=	2831	;
conv3_kernel[0][1][1][3]=	281	;
conv3_kernel[0][1][1][4]=	-283	;
conv3_kernel[0][1][2][0]=	-6147	;
conv3_kernel[0][1][2][1]=	-547	;
conv3_kernel[0][1][2][2]=	3500	;
conv3_kernel[0][1][2][3]=	3203	;
conv3_kernel[0][1][2][4]=	-6028	;
conv3_kernel[0][1][3][0]=	6819	;
conv3_kernel[0][1][3][1]=	390	;
conv3_kernel[0][1][3][2]=	-383	;
conv3_kernel[0][1][3][3]=	-2143	;
conv3_kernel[0][1][3][4]=	3149	;
conv3_kernel[0][1][4][0]=	10524	;
conv3_kernel[0][1][4][1]=	-2552	;
conv3_kernel[0][1][4][2]=	473	;
conv3_kernel[0][1][4][3]=	1670	;
conv3_kernel[0][1][4][4]=	6385	;
conv3_kernel[1][0][0][0]=	4740	;
conv3_kernel[1][0][0][1]=	2421	;
conv3_kernel[1][0][0][2]=	-680	;
conv3_kernel[1][0][0][3]=	-1782	;
conv3_kernel[1][0][0][4]=	-10590	;
conv3_kernel[1][0][1][0]=	1591	;
conv3_kernel[1][0][1][1]=	1540	;
conv3_kernel[1][0][1][2]=	-1481	;
conv3_kernel[1][0][1][3]=	-489	;
conv3_kernel[1][0][1][4]=	-10351	;
conv3_kernel[1][0][2][0]=	-6423	;
conv3_kernel[1][0][2][1]=	-1419	;
conv3_kernel[1][0][2][2]=	-87	;
conv3_kernel[1][0][2][3]=	313	;
conv3_kernel[1][0][2][4]=	6857	;
conv3_kernel[1][0][3][0]=	-3169	;
conv3_kernel[1][0][3][1]=	3640	;
conv3_kernel[1][0][3][2]=	5005	;
conv3_kernel[1][0][3][3]=	-131	;
conv3_kernel[1][0][3][4]=	5296	;
conv3_kernel[1][0][4][0]=	5019	;
conv3_kernel[1][0][4][1]=	4779	;
conv3_kernel[1][0][4][2]=	-1042	;
conv3_kernel[1][0][4][3]=	-1350	;
conv3_kernel[1][0][4][4]=	-623	;
conv3_kernel[1][1][0][0]=	-3313	;
conv3_kernel[1][1][0][1]=	-3189	;
conv3_kernel[1][1][0][2]=	-1487	;
conv3_kernel[1][1][0][3]=	-843	;
conv3_kernel[1][1][0][4]=	2935	;
conv3_kernel[1][1][1][0]=	2711	;
conv3_kernel[1][1][1][1]=	-749	;
conv3_kernel[1][1][1][2]=	-2549	;
conv3_kernel[1][1][1][3]=	3076	;
conv3_kernel[1][1][1][4]=	1725	;
conv3_kernel[1][1][2][0]=	3231	;
conv3_kernel[1][1][2][1]=	904	;
conv3_kernel[1][1][2][2]=	-1828	;
conv3_kernel[1][1][2][3]=	4389	;
conv3_kernel[1][1][2][4]=	-2104	;
conv3_kernel[1][1][3][0]=	-4469	;
conv3_kernel[1][1][3][1]=	3354	;
conv3_kernel[1][1][3][2]=	-1590	;
conv3_kernel[1][1][3][3]=	-709	;
conv3_kernel[1][1][3][4]=	2107	;
conv3_kernel[1][1][4][0]=	-11487	;
conv3_kernel[1][1][4][1]=	2667	;
conv3_kernel[1][1][4][2]=	1816	;
conv3_kernel[1][1][4][3]=	5558	;
conv3_kernel[1][1][4][4]=	5054	;
conv3_kernel[2][0][0][0]=	3831	;
conv3_kernel[2][0][0][1]=	5347	;
conv3_kernel[2][0][0][2]=	-2045	;
conv3_kernel[2][0][0][3]=	2241	;
conv3_kernel[2][0][0][4]=	-4713	;
conv3_kernel[2][0][1][0]=	-2017	;
conv3_kernel[2][0][1][1]=	1781	;
conv3_kernel[2][0][1][2]=	1229	;
conv3_kernel[2][0][1][3]=	-363	;
conv3_kernel[2][0][1][4]=	-5531	;
conv3_kernel[2][0][2][0]=	951	;
conv3_kernel[2][0][2][1]=	957	;
conv3_kernel[2][0][2][2]=	-1437	;
conv3_kernel[2][0][2][3]=	7563	;
conv3_kernel[2][0][2][4]=	4443	;
conv3_kernel[2][0][3][0]=	1160	;
conv3_kernel[2][0][3][1]=	-244	;
conv3_kernel[2][0][3][2]=	252	;
conv3_kernel[2][0][3][3]=	7538	;
conv3_kernel[2][0][3][4]=	2230	;
conv3_kernel[2][0][4][0]=	-824	;
conv3_kernel[2][0][4][1]=	-2753	;
conv3_kernel[2][0][4][2]=	-3827	;
conv3_kernel[2][0][4][3]=	-472	;
conv3_kernel[2][0][4][4]=	1916	;
conv3_kernel[2][1][0][0]=	-198	;
conv3_kernel[2][1][0][1]=	12	;
conv3_kernel[2][1][0][2]=	1003	;
conv3_kernel[2][1][0][3]=	-32	;
conv3_kernel[2][1][0][4]=	1901	;
conv3_kernel[2][1][1][0]=	3689	;
conv3_kernel[2][1][1][1]=	1291	;
conv3_kernel[2][1][1][2]=	1430	;
conv3_kernel[2][1][1][3]=	3692	;
conv3_kernel[2][1][1][4]=	1233	;
conv3_kernel[2][1][2][0]=	-3128	;
conv3_kernel[2][1][2][1]=	-770	;
conv3_kernel[2][1][2][2]=	1191	;
conv3_kernel[2][1][2][3]=	6030	;
conv3_kernel[2][1][2][4]=	-5743	;
conv3_kernel[2][1][3][0]=	-900	;
conv3_kernel[2][1][3][1]=	849	;
conv3_kernel[2][1][3][2]=	1952	;
conv3_kernel[2][1][3][3]=	-3841	;
conv3_kernel[2][1][3][4]=	-4443	;
conv3_kernel[2][1][4][0]=	3210	;
conv3_kernel[2][1][4][1]=	-2036	;
conv3_kernel[2][1][4][2]=	-4338	;
conv3_kernel[2][1][4][3]=	-865	;
conv3_kernel[2][1][4][4]=	-152	;
conv3_kernel[3][0][0][0]=	1286	;
conv3_kernel[3][0][0][1]=	-2043	;
conv3_kernel[3][0][0][2]=	1625	;
conv3_kernel[3][0][0][3]=	-1714	;
conv3_kernel[3][0][0][4]=	-2583	;
conv3_kernel[3][0][1][0]=	2783	;
conv3_kernel[3][0][1][1]=	-1434	;
conv3_kernel[3][0][1][2]=	-59	;
conv3_kernel[3][0][1][3]=	152	;
conv3_kernel[3][0][1][4]=	4407	;
conv3_kernel[3][0][2][0]=	-93	;
conv3_kernel[3][0][2][1]=	-4078	;
conv3_kernel[3][0][2][2]=	72	;
conv3_kernel[3][0][2][3]=	3275	;
conv3_kernel[3][0][2][4]=	2219	;
conv3_kernel[3][0][3][0]=	-2502	;
conv3_kernel[3][0][3][1]=	-1172	;
conv3_kernel[3][0][3][2]=	2109	;
conv3_kernel[3][0][3][3]=	-7488	;
conv3_kernel[3][0][3][4]=	-1185	;
conv3_kernel[3][0][4][0]=	4191	;
conv3_kernel[3][0][4][1]=	2480	;
conv3_kernel[3][0][4][2]=	3756	;
conv3_kernel[3][0][4][3]=	-848	;
conv3_kernel[3][0][4][4]=	-4081	;
conv3_kernel[3][1][0][0]=	2132	;
conv3_kernel[3][1][0][1]=	1029	;
conv3_kernel[3][1][0][2]=	1067	;
conv3_kernel[3][1][0][3]=	-5153	;
conv3_kernel[3][1][0][4]=	2197	;
conv3_kernel[3][1][1][0]=	-1679	;
conv3_kernel[3][1][1][1]=	232	;
conv3_kernel[3][1][1][2]=	2015	;
conv3_kernel[3][1][1][3]=	1588	;
conv3_kernel[3][1][1][4]=	-828	;
conv3_kernel[3][1][2][0]=	-2024	;
conv3_kernel[3][1][2][1]=	8	;
conv3_kernel[3][1][2][2]=	7592	;
conv3_kernel[3][1][2][3]=	5420	;
conv3_kernel[3][1][2][4]=	3737	;
conv3_kernel[3][1][3][0]=	8432	;
conv3_kernel[3][1][3][1]=	-1032	;
conv3_kernel[3][1][3][2]=	-1190	;
conv3_kernel[3][1][3][3]=	2413	;
conv3_kernel[3][1][3][4]=	6988	;
conv3_kernel[3][1][4][0]=	-15493	;
conv3_kernel[3][1][4][1]=	-1687	;
conv3_kernel[3][1][4][2]=	1464	;
conv3_kernel[3][1][4][3]=	1593	;
conv3_kernel[3][1][4][4]=	-1473	;
conv3_kernel[4][0][0][0]=	-974	;
conv3_kernel[4][0][0][1]=	4120	;
conv3_kernel[4][0][0][2]=	6341	;
conv3_kernel[4][0][0][3]=	9967	;
conv3_kernel[4][0][0][4]=	6357	;
conv3_kernel[4][0][1][0]=	1220	;
conv3_kernel[4][0][1][1]=	473	;
conv3_kernel[4][0][1][2]=	699	;
conv3_kernel[4][0][1][3]=	1439	;
conv3_kernel[4][0][1][4]=	3087	;
conv3_kernel[4][0][2][0]=	-3227	;
conv3_kernel[4][0][2][1]=	-978	;
conv3_kernel[4][0][2][2]=	2841	;
conv3_kernel[4][0][2][3]=	-4558	;
conv3_kernel[4][0][2][4]=	-5782	;
conv3_kernel[4][0][3][0]=	-1231	;
conv3_kernel[4][0][3][1]=	181	;
conv3_kernel[4][0][3][2]=	4702	;
conv3_kernel[4][0][3][3]=	-3039	;
conv3_kernel[4][0][3][4]=	-136	;
conv3_kernel[4][0][4][0]=	1094	;
conv3_kernel[4][0][4][1]=	-1426	;
conv3_kernel[4][0][4][2]=	2519	;
conv3_kernel[4][0][4][3]=	703	;
conv3_kernel[4][0][4][4]=	-3684	;
conv3_kernel[4][1][0][0]=	2762	;
conv3_kernel[4][1][0][1]=	-1952	;
conv3_kernel[4][1][0][2]=	-4382	;
conv3_kernel[4][1][0][3]=	-9609	;
conv3_kernel[4][1][0][4]=	-2240	;
conv3_kernel[4][1][1][0]=	-2695	;
conv3_kernel[4][1][1][1]=	-1717	;
conv3_kernel[4][1][1][2]=	-853	;
conv3_kernel[4][1][1][3]=	1790	;
conv3_kernel[4][1][1][4]=	9329	;
conv3_kernel[4][1][2][0]=	-4747	;
conv3_kernel[4][1][2][1]=	752	;
conv3_kernel[4][1][2][2]=	3924	;
conv3_kernel[4][1][2][3]=	6416	;
conv3_kernel[4][1][2][4]=	6147	;
conv3_kernel[4][1][3][0]=	-446	;
conv3_kernel[4][1][3][1]=	4227	;
conv3_kernel[4][1][3][2]=	607	;
conv3_kernel[4][1][3][3]=	2241	;
conv3_kernel[4][1][3][4]=	-1254	;
conv3_kernel[4][1][4][0]=	-4419	;
conv3_kernel[4][1][4][1]=	2932	;
conv3_kernel[4][1][4][2]=	1571	;
conv3_kernel[4][1][4][3]=	3282	;
conv3_kernel[4][1][4][4]=	-335	;
conv3_kernel[5][0][0][0]=	9875	;
conv3_kernel[5][0][0][1]=	4267	;
conv3_kernel[5][0][0][2]=	2953	;
conv3_kernel[5][0][0][3]=	-2185	;
conv3_kernel[5][0][0][4]=	-4306	;
conv3_kernel[5][0][1][0]=	5698	;
conv3_kernel[5][0][1][1]=	1489	;
conv3_kernel[5][0][1][2]=	466	;
conv3_kernel[5][0][1][3]=	-428	;
conv3_kernel[5][0][1][4]=	1063	;
conv3_kernel[5][0][2][0]=	1899	;
conv3_kernel[5][0][2][1]=	-788	;
conv3_kernel[5][0][2][2]=	-1123	;
conv3_kernel[5][0][2][3]=	325	;
conv3_kernel[5][0][2][4]=	-2858	;
conv3_kernel[5][0][3][0]=	-3	;
conv3_kernel[5][0][3][1]=	1656	;
conv3_kernel[5][0][3][2]=	-1176	;
conv3_kernel[5][0][3][3]=	-367	;
conv3_kernel[5][0][3][4]=	-251	;
conv3_kernel[5][0][4][0]=	410	;
conv3_kernel[5][0][4][1]=	-2999	;
conv3_kernel[5][0][4][2]=	-2942	;
conv3_kernel[5][0][4][3]=	1074	;
conv3_kernel[5][0][4][4]=	-4413	;
conv3_kernel[5][1][0][0]=	-5603	;
conv3_kernel[5][1][0][1]=	652	;
conv3_kernel[5][1][0][2]=	2063	;
conv3_kernel[5][1][0][3]=	-362	;
conv3_kernel[5][1][0][4]=	754	;
conv3_kernel[5][1][1][0]=	-2285	;
conv3_kernel[5][1][1][1]=	3934	;
conv3_kernel[5][1][1][2]=	1479	;
conv3_kernel[5][1][1][3]=	2640	;
conv3_kernel[5][1][1][4]=	1145	;
conv3_kernel[5][1][2][0]=	7751	;
conv3_kernel[5][1][2][1]=	-909	;
conv3_kernel[5][1][2][2]=	199	;
conv3_kernel[5][1][2][3]=	2351	;
conv3_kernel[5][1][2][4]=	4779	;
conv3_kernel[5][1][3][0]=	12350	;
conv3_kernel[5][1][3][1]=	1497	;
conv3_kernel[5][1][3][2]=	-1655	;
conv3_kernel[5][1][3][3]=	3076	;
conv3_kernel[5][1][3][4]=	1266	;
conv3_kernel[5][1][4][0]=	10776	;
conv3_kernel[5][1][4][1]=	3231	;
conv3_kernel[5][1][4][2]=	2458	;
conv3_kernel[5][1][4][3]=	259	;
conv3_kernel[5][1][4][4]=	-2695	;
conv3_kernel[6][0][0][0]=	-1462	;
conv3_kernel[6][0][0][1]=	-5954	;
conv3_kernel[6][0][0][2]=	-3058	;
conv3_kernel[6][0][0][3]=	726	;
conv3_kernel[6][0][0][4]=	4434	;
conv3_kernel[6][0][1][0]=	-1975	;
conv3_kernel[6][0][1][1]=	2207	;
conv3_kernel[6][0][1][2]=	1151	;
conv3_kernel[6][0][1][3]=	1140	;
conv3_kernel[6][0][1][4]=	2988	;
conv3_kernel[6][0][2][0]=	2219	;
conv3_kernel[6][0][2][1]=	-234	;
conv3_kernel[6][0][2][2]=	-1752	;
conv3_kernel[6][0][2][3]=	7479	;
conv3_kernel[6][0][2][4]=	2337	;
conv3_kernel[6][0][3][0]=	-1058	;
conv3_kernel[6][0][3][1]=	2355	;
conv3_kernel[6][0][3][2]=	-809	;
conv3_kernel[6][0][3][3]=	3078	;
conv3_kernel[6][0][3][4]=	4828	;
conv3_kernel[6][0][4][0]=	3864	;
conv3_kernel[6][0][4][1]=	-1445	;
conv3_kernel[6][0][4][2]=	-61	;
conv3_kernel[6][0][4][3]=	1123	;
conv3_kernel[6][0][4][4]=	-1216	;
conv3_kernel[6][1][0][0]=	5573	;
conv3_kernel[6][1][0][1]=	968	;
conv3_kernel[6][1][0][2]=	-3960	;
conv3_kernel[6][1][0][3]=	-9163	;
conv3_kernel[6][1][0][4]=	-4700	;
conv3_kernel[6][1][1][0]=	-2613	;
conv3_kernel[6][1][1][1]=	243	;
conv3_kernel[6][1][1][2]=	-816	;
conv3_kernel[6][1][1][3]=	-1350	;
conv3_kernel[6][1][1][4]=	-1175	;
conv3_kernel[6][1][2][0]=	5049	;
conv3_kernel[6][1][2][1]=	1710	;
conv3_kernel[6][1][2][2]=	2245	;
conv3_kernel[6][1][2][3]=	8683	;
conv3_kernel[6][1][2][4]=	1270	;
conv3_kernel[6][1][3][0]=	5745	;
conv3_kernel[6][1][3][1]=	1933	;
conv3_kernel[6][1][3][2]=	1203	;
conv3_kernel[6][1][3][3]=	2864	;
conv3_kernel[6][1][3][4]=	6220	;
conv3_kernel[6][1][4][0]=	-3976	;
conv3_kernel[6][1][4][1]=	-1968	;
conv3_kernel[6][1][4][2]=	-1469	;
conv3_kernel[6][1][4][3]=	-5043	;
conv3_kernel[6][1][4][4]=	2835	;
conv3_kernel[7][0][0][0]=	-1931	;
conv3_kernel[7][0][0][1]=	-66	;
conv3_kernel[7][0][0][2]=	-5311	;
conv3_kernel[7][0][0][3]=	-2760	;
conv3_kernel[7][0][0][4]=	-506	;
conv3_kernel[7][0][1][0]=	-9080	;
conv3_kernel[7][0][1][1]=	559	;
conv3_kernel[7][0][1][2]=	2316	;
conv3_kernel[7][0][1][3]=	1156	;
conv3_kernel[7][0][1][4]=	516	;
conv3_kernel[7][0][2][0]=	1648	;
conv3_kernel[7][0][2][1]=	1592	;
conv3_kernel[7][0][2][2]=	1098	;
conv3_kernel[7][0][2][3]=	905	;
conv3_kernel[7][0][2][4]=	2108	;
conv3_kernel[7][0][3][0]=	3147	;
conv3_kernel[7][0][3][1]=	365	;
conv3_kernel[7][0][3][2]=	-283	;
conv3_kernel[7][0][3][3]=	-2956	;
conv3_kernel[7][0][3][4]=	-7987	;
conv3_kernel[7][0][4][0]=	-300	;
conv3_kernel[7][0][4][1]=	305	;
conv3_kernel[7][0][4][2]=	-1848	;
conv3_kernel[7][0][4][3]=	825	;
conv3_kernel[7][0][4][4]=	4263	;
conv3_kernel[7][1][0][0]=	1237	;
conv3_kernel[7][1][0][1]=	5158	;
conv3_kernel[7][1][0][2]=	646	;
conv3_kernel[7][1][0][3]=	220	;
conv3_kernel[7][1][0][4]=	4460	;
conv3_kernel[7][1][1][0]=	5007	;
conv3_kernel[7][1][1][1]=	616	;
conv3_kernel[7][1][1][2]=	1085	;
conv3_kernel[7][1][1][3]=	1121	;
conv3_kernel[7][1][1][4]=	1875	;
conv3_kernel[7][1][2][0]=	-4787	;
conv3_kernel[7][1][2][1]=	-3465	;
conv3_kernel[7][1][2][2]=	4363	;
conv3_kernel[7][1][2][3]=	7133	;
conv3_kernel[7][1][2][4]=	-823	;
conv3_kernel[7][1][3][0]=	-2955	;
conv3_kernel[7][1][3][1]=	3041	;
conv3_kernel[7][1][3][2]=	4530	;
conv3_kernel[7][1][3][3]=	2750	;
conv3_kernel[7][1][3][4]=	-5431	;
conv3_kernel[7][1][4][0]=	4704	;
conv3_kernel[7][1][4][1]=	2587	;
conv3_kernel[7][1][4][2]=	3467	;
conv3_kernel[7][1][4][3]=	-1308	;
conv3_kernel[7][1][4][4]=	-8905	;
conv3_kernel[8][0][0][0]=	-9776	;
conv3_kernel[8][0][0][1]=	-3763	;
conv3_kernel[8][0][0][2]=	1900	;
conv3_kernel[8][0][0][3]=	-426	;
conv3_kernel[8][0][0][4]=	2838	;
conv3_kernel[8][0][1][0]=	-14842	;
conv3_kernel[8][0][1][1]=	317	;
conv3_kernel[8][0][1][2]=	273	;
conv3_kernel[8][0][1][3]=	613	;
conv3_kernel[8][0][1][4]=	-1007	;
conv3_kernel[8][0][2][0]=	2856	;
conv3_kernel[8][0][2][1]=	-2307	;
conv3_kernel[8][0][2][2]=	2039	;
conv3_kernel[8][0][2][3]=	1652	;
conv3_kernel[8][0][2][4]=	5176	;
conv3_kernel[8][0][3][0]=	-296	;
conv3_kernel[8][0][3][1]=	-384	;
conv3_kernel[8][0][3][2]=	1238	;
conv3_kernel[8][0][3][3]=	-1976	;
conv3_kernel[8][0][3][4]=	-360	;
conv3_kernel[8][0][4][0]=	2266	;
conv3_kernel[8][0][4][1]=	894	;
conv3_kernel[8][0][4][2]=	-276	;
conv3_kernel[8][0][4][3]=	994	;
conv3_kernel[8][0][4][4]=	-639	;
conv3_kernel[8][1][0][0]=	7340	;
conv3_kernel[8][1][0][1]=	5169	;
conv3_kernel[8][1][0][2]=	398	;
conv3_kernel[8][1][0][3]=	-822	;
conv3_kernel[8][1][0][4]=	3897	;
conv3_kernel[8][1][1][0]=	3251	;
conv3_kernel[8][1][1][1]=	834	;
conv3_kernel[8][1][1][2]=	1308	;
conv3_kernel[8][1][1][3]=	3487	;
conv3_kernel[8][1][1][4]=	4021	;
conv3_kernel[8][1][2][0]=	753	;
conv3_kernel[8][1][2][1]=	-4231	;
conv3_kernel[8][1][2][2]=	-5108	;
conv3_kernel[8][1][2][3]=	-2006	;
conv3_kernel[8][1][2][4]=	-4125	;
conv3_kernel[8][1][3][0]=	-2236	;
conv3_kernel[8][1][3][1]=	-1804	;
conv3_kernel[8][1][3][2]=	-2033	;
conv3_kernel[8][1][3][3]=	-43	;
conv3_kernel[8][1][3][4]=	-3445	;
conv3_kernel[8][1][4][0]=	-9703	;
conv3_kernel[8][1][4][1]=	1211	;
conv3_kernel[8][1][4][2]=	1140	;
conv3_kernel[8][1][4][3]=	1345	;
conv3_kernel[8][1][4][4]=	-7669	;
conv3_kernel[9][0][0][0]=	5466	;
conv3_kernel[9][0][0][1]=	-3611	;
conv3_kernel[9][0][0][2]=	-3640	;
conv3_kernel[9][0][0][3]=	-6320	;
conv3_kernel[9][0][0][4]=	-3012	;
conv3_kernel[9][0][1][0]=	5214	;
conv3_kernel[9][0][1][1]=	-2271	;
conv3_kernel[9][0][1][2]=	2164	;
conv3_kernel[9][0][1][3]=	2329	;
conv3_kernel[9][0][1][4]=	1095	;
conv3_kernel[9][0][2][0]=	-404	;
conv3_kernel[9][0][2][1]=	-1823	;
conv3_kernel[9][0][2][2]=	8974	;
conv3_kernel[9][0][2][3]=	5216	;
conv3_kernel[9][0][2][4]=	53	;
conv3_kernel[9][0][3][0]=	-2398	;
conv3_kernel[9][0][3][1]=	-2000	;
conv3_kernel[9][0][3][2]=	5404	;
conv3_kernel[9][0][3][3]=	-3861	;
conv3_kernel[9][0][3][4]=	132	;
conv3_kernel[9][0][4][0]=	460	;
conv3_kernel[9][0][4][1]=	-4874	;
conv3_kernel[9][0][4][2]=	5580	;
conv3_kernel[9][0][4][3]=	3040	;
conv3_kernel[9][0][4][4]=	-2862	;
conv3_kernel[9][1][0][0]=	-933	;
conv3_kernel[9][1][0][1]=	1661	;
conv3_kernel[9][1][0][2]=	5667	;
conv3_kernel[9][1][0][3]=	-4670	;
conv3_kernel[9][1][0][4]=	-1087	;
conv3_kernel[9][1][1][0]=	-589	;
conv3_kernel[9][1][1][1]=	-1588	;
conv3_kernel[9][1][1][2]=	1456	;
conv3_kernel[9][1][1][3]=	-3259	;
conv3_kernel[9][1][1][4]=	-4431	;
conv3_kernel[9][1][2][0]=	-313	;
conv3_kernel[9][1][2][1]=	-1521	;
conv3_kernel[9][1][2][2]=	3676	;
conv3_kernel[9][1][2][3]=	-420	;
conv3_kernel[9][1][2][4]=	-153	;
conv3_kernel[9][1][3][0]=	2170	;
conv3_kernel[9][1][3][1]=	863	;
conv3_kernel[9][1][3][2]=	544	;
conv3_kernel[9][1][3][3]=	483	;
conv3_kernel[9][1][3][4]=	354	;
conv3_kernel[9][1][4][0]=	1832	;
conv3_kernel[9][1][4][1]=	3393	;
conv3_kernel[9][1][4][2]=	143	;
conv3_kernel[9][1][4][3]=	-455	;
conv3_kernel[9][1][4][4]=	-1689	;
connect_matrix [0][0]=	-5549	;
connect_matrix [0][1]=	6296	;
connect_matrix [0][2]=	-863	;
connect_matrix [0][3]=	-4980	;
connect_matrix [0][4]=	835	;
connect_matrix [0][5]=	-988	;
connect_matrix [0][6]=	-341	;
connect_matrix [0][7]=	-231	;
connect_matrix [0][8]=	3243	;
connect_matrix [0][9]=	-3070	;
connect_matrix [1][0]=	6852	;
connect_matrix [1][1]=	-2251	;
connect_matrix [1][2]=	-6471	;
connect_matrix [1][3]=	-5020	;
connect_matrix [1][4]=	-30	;
connect_matrix [1][5]=	2448	;
connect_matrix [1][6]=	2564	;
connect_matrix [1][7]=	-12052	;
connect_matrix [1][8]=	6356	;
connect_matrix [1][9]=	9423	;
connect_matrix [2][0]=	2618	;
connect_matrix [2][1]=	5434	;
connect_matrix [2][2]=	-241	;
connect_matrix [2][3]=	2375	;
connect_matrix [2][4]=	-5801	;
connect_matrix [2][5]=	3131	;
connect_matrix [2][6]=	732	;
connect_matrix [2][7]=	-2819	;
connect_matrix [2][8]=	-7247	;
connect_matrix [2][9]=	-336	;
connect_matrix [3][0]=	-1747	;
connect_matrix [3][1]=	-197	;
connect_matrix [3][2]=	-4129	;
connect_matrix [3][3]=	-68	;
connect_matrix [3][4]=	-1102	;
connect_matrix [3][5]=	6075	;
connect_matrix [3][6]=	-1689	;
connect_matrix [3][7]=	2787	;
connect_matrix [3][8]=	-5818	;
connect_matrix [3][9]=	2854	;
connect_matrix [4][0]=	-29	;
connect_matrix [4][1]=	-2343	;
connect_matrix [4][2]=	-702	;
connect_matrix [4][3]=	-2113	;
connect_matrix [4][4]=	-4308	;
connect_matrix [4][5]=	-5942	;
connect_matrix [4][6]=	8167	;
connect_matrix [4][7]=	3606	;
connect_matrix [4][8]=	-2518	;
connect_matrix [4][9]=	2918	;
connect_matrix [5][0]=	2274	;
connect_matrix [5][1]=	-4095	;
connect_matrix [5][2]=	-4361	;
connect_matrix [5][3]=	-1600	;
connect_matrix [5][4]=	5423	;
connect_matrix [5][5]=	3144	;
connect_matrix [5][6]=	-935	;
connect_matrix [5][7]=	2530	;
connect_matrix [5][8]=	-810	;
connect_matrix [5][9]=	-4821	;
connect_matrix [6][0]=	-6693	;
connect_matrix [6][1]=	3317	;
connect_matrix [6][2]=	2632	;
connect_matrix [6][3]=	1190	;
connect_matrix [6][4]=	7894	;
connect_matrix [6][5]=	-11649	;
connect_matrix [6][6]=	1658	;
connect_matrix [6][7]=	-1742	;
connect_matrix [6][8]=	-1846	;
connect_matrix [6][9]=	-1999	;
connect_matrix [7][0]=	-4040	;
connect_matrix [7][1]=	-5540	;
connect_matrix [7][2]=	6922	;
connect_matrix [7][3]=	2518	;
connect_matrix [7][4]=	-625	;
connect_matrix [7][5]=	3608	;
connect_matrix [7][6]=	-45	;
connect_matrix [7][7]=	-4983	;
connect_matrix [7][8]=	3509	;
connect_matrix [7][9]=	2141	;
connect_matrix [8][0]=	884	;
connect_matrix [8][1]=	-258	;
connect_matrix [8][2]=	305	;
connect_matrix [8][3]=	7368	;
connect_matrix [8][4]=	-1753	;
connect_matrix [8][5]=	-1196	;
connect_matrix [8][6]=	-3660	;
connect_matrix [8][7]=	1489	;
connect_matrix [8][8]=	1440	;
connect_matrix [8][9]=	-1175	;
connect_matrix [9][0]=	3438	;
connect_matrix [9][1]=	-892	;
connect_matrix [9][2]=	4805	;
connect_matrix [9][3]=	-2545	;
connect_matrix [9][4]=	-1441	;
connect_matrix [9][5]=	-2977	;
connect_matrix [9][6]=	-4518	;
connect_matrix [9][7]=	5422	;
connect_matrix [9][8]=	-4027	;
connect_matrix [9][9]=	2192	;
end
endmodule